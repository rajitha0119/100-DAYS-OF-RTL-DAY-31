`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 24.08.2023 22:18:15
// Design Name: 
// Module Name: pipo
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module d_ff(input clk, input d,output reg q);
always@(negedge clk or d)
begin
q<=d;
end
endmodule

module pipo(
    input clk,
    input [3:0]d,
    output reg [3:0]q
    );
    d_ff DFF1(clk,d[3],q[3]);
    d_ff DFF2(clk,d[2],q[2]);
    d_ff DFF3(clk,d[1],q[1]);
    d_ff DFF4(clk.d[0],q[0]);
endmodule
